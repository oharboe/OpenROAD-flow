module ibex_cs_registers (
	clk_i,
	rst_ni,
	hart_id_i,
	priv_mode_id_o,
	priv_mode_if_o,
	priv_mode_lsu_o,
	csr_mstatus_tw_o,
	csr_mtvec_o,
	csr_mtvec_init_i,
	boot_addr_i,
	csr_access_i,
	csr_addr_i,
	csr_wdata_i,
	csr_op_i,
	csr_rdata_o,
	irq_software_i,
	irq_timer_i,
	irq_external_i,
	irq_fast_i,
	irq_pending_o,
	csr_msip_o,
	csr_mtip_o,
	csr_meip_o,
	csr_mfip_o,
	csr_mstatus_mie_o,
	csr_mepc_o,
	csr_pmp_cfg_o,
	csr_pmp_addr_o,
	debug_mode_i,
	debug_cause_i,
	debug_csr_save_i,
	csr_depc_o,
	debug_single_step_o,
	debug_ebreakm_o,
	debug_ebreaku_o,
	pc_if_i,
	pc_id_i,
	csr_save_if_i,
	csr_save_id_i,
	csr_restore_mret_i,
	csr_save_cause_i,
	csr_mcause_i,
	csr_mtval_i,
	illegal_csr_insn_o,
	instr_new_id_i,
	instr_ret_i,
	instr_ret_compressed_i,
	imiss_i,
	pc_set_i,
	jump_i,
	branch_i,
	branch_taken_i,
	mem_load_i,
	mem_store_i,
	lsu_busy_i
);
	parameter [31:0] MHPMCounterNum = 8;
	parameter [31:0] MHPMCounterWidth = 40;
	parameter PMPEnable = 0;
	parameter [31:0] PMPGranularity = 0;
	parameter [31:0] PMPNumRegions = 4;
	parameter RV32E = 0;
	parameter RV32M = 0;
	input wire clk_i;
	input wire rst_ni;
	input wire [31:0] hart_id_i;
	output wire [1:0] priv_mode_id_o;
	output wire [1:0] priv_mode_if_o;
	output wire [1:0] priv_mode_lsu_o;
	output wire csr_mstatus_tw_o;
	output wire [31:0] csr_mtvec_o;
	input wire csr_mtvec_init_i;
	input wire [31:0] boot_addr_i;
	input wire csr_access_i;
	input wire [11:0] csr_addr_i;
	input wire [31:0] csr_wdata_i;
	input wire [1:0] csr_op_i;
	output wire [31:0] csr_rdata_o;
	input wire irq_software_i;
	input wire irq_timer_i;
	input wire irq_external_i;
	input wire [14:0] irq_fast_i;
	output wire irq_pending_o;
	output wire csr_msip_o;
	output wire csr_mtip_o;
	output wire csr_meip_o;
	output wire [14:0] csr_mfip_o;
	output wire csr_mstatus_mie_o;
	output wire [31:0] csr_mepc_o;
	output wire [((0 >= (PMPNumRegions - 1)) ? ((((0 >= (PMPNumRegions - 1)) ? (2 - PMPNumRegions) : PMPNumRegions) * 6) + (((PMPNumRegions - 1) * 6) - 1)) : (((((PMPNumRegions - 1) >= 0) ? PMPNumRegions : (2 - PMPNumRegions)) * 6) + -1)):((0 >= (PMPNumRegions - 1)) ? ((PMPNumRegions - 1) * 6) : 0)] csr_pmp_cfg_o;
	output wire [((0 >= (PMPNumRegions - 1)) ? ((((0 >= (PMPNumRegions - 1)) ? (2 - PMPNumRegions) : PMPNumRegions) * 34) + (((PMPNumRegions - 1) * 34) - 1)) : (((((PMPNumRegions - 1) >= 0) ? PMPNumRegions : (2 - PMPNumRegions)) * 34) + -1)):((0 >= (PMPNumRegions - 1)) ? ((PMPNumRegions - 1) * 34) : 0)] csr_pmp_addr_o;
	input wire debug_mode_i;
	input wire [2:0] debug_cause_i;
	input wire debug_csr_save_i;
	output wire [31:0] csr_depc_o;
	output wire debug_single_step_o;
	output wire debug_ebreakm_o;
	output wire debug_ebreaku_o;
	input wire [31:0] pc_if_i;
	input wire [31:0] pc_id_i;
	input wire csr_save_if_i;
	input wire csr_save_id_i;
	input wire csr_restore_mret_i;
	input wire csr_save_cause_i;
	input wire [5:0] csr_mcause_i;
	input wire [31:0] csr_mtval_i;
	output wire illegal_csr_insn_o;
	input wire instr_new_id_i;
	input wire instr_ret_i;
	input wire instr_ret_compressed_i;
	input wire imiss_i;
	input wire pc_set_i;
	input wire jump_i;
	input wire branch_i;
	input wire branch_taken_i;
	input wire mem_load_i;
	input wire mem_store_i;
	input wire lsu_busy_i;
	parameter [31:0] PMP_MAX_REGIONS = 16;
	parameter [31:0] PMP_CFG_W = 8;
	parameter [31:0] PMP_I = 0;
	parameter [31:0] PMP_D = 1;
	parameter [11:0] CSR_OFF_PMP_CFG = 12'h3A0;
	parameter [11:0] CSR_OFF_PMP_ADDR = 12'h3B0;
	parameter [11:0] CSR_OFF_MCOUNTER_SETUP = 12'h320;
	parameter [11:0] CSR_OFF_MCOUNTER = 12'hB00;
	parameter [11:0] CSR_OFF_MCOUNTERH = 12'hB80;
	parameter [11:0] CSR_MASK_MCOUNTER = 12'hFE0;
	parameter [31:0] CSR_MSTATUS_MIE_BIT = 3;
	parameter [31:0] CSR_MSTATUS_MPIE_BIT = 7;
	parameter [31:0] CSR_MSTATUS_MPP_BIT_LOW = 11;
	parameter [31:0] CSR_MSTATUS_MPP_BIT_HIGH = 12;
	parameter [31:0] CSR_MSTATUS_MPRV_BIT = 17;
	parameter [31:0] CSR_MSTATUS_TW_BIT = 21;
	parameter [31:0] CSR_MSIX_BIT = 3;
	parameter [31:0] CSR_MTIX_BIT = 7;
	parameter [31:0] CSR_MEIX_BIT = 11;
	parameter [31:0] CSR_MFIX_BIT_LOW = 16;
	parameter [31:0] CSR_MFIX_BIT_HIGH = 30;
	localparam [0:0] IMM_A_Z = 0;
	localparam [0:0] OP_B_REG_B = 0;
	localparam [1:0] CSR_OP_READ = 0;
	localparam [1:0] EXC_PC_EXC = 0;
	localparam [1:0] MD_OP_MULL = 0;
	localparam [1:0] OP_A_REG_A = 0;
	localparam [1:0] RF_WD_LSU = 0;
	localparam [2:0] IMM_B_I = 0;
	localparam [2:0] PC_BOOT = 0;
	localparam [4:0] ALU_ADD = 0;
	localparam [0:0] IMM_A_ZERO = 1;
	localparam [0:0] OP_B_IMM = 1;
	localparam [1:0] CSR_OP_WRITE = 1;
	localparam [1:0] EXC_PC_IRQ = 1;
	localparam [1:0] MD_OP_MULH = 1;
	localparam [1:0] OP_A_FWD = 1;
	localparam [1:0] RF_WD_EX = 1;
	localparam [2:0] IMM_B_S = 1;
	localparam [2:0] PC_JUMP = 1;
	localparam [4:0] ALU_SUB = 1;
	localparam [4:0] ALU_LE = 10;
	localparam [4:0] ALU_LEU = 11;
	localparam [4:0] ALU_GT = 12;
	localparam [11:0] CSR_MSTATUS = 12'h300;
	localparam [11:0] CSR_MISA = 12'h301;
	localparam [11:0] CSR_MIE = 12'h304;
	localparam [11:0] CSR_MTVEC = 12'h305;
	localparam [11:0] CSR_MCOUNTINHIBIT = 12'h320;
	localparam [11:0] CSR_MSCRATCH = 12'h340;
	localparam [11:0] CSR_MEPC = 12'h341;
	localparam [11:0] CSR_MCAUSE = 12'h342;
	localparam [11:0] CSR_MTVAL = 12'h343;
	localparam [11:0] CSR_MIP = 12'h344;
	localparam [11:0] CSR_PMPCFG0 = 12'h3A0;
	localparam [11:0] CSR_PMPCFG1 = 12'h3A1;
	localparam [11:0] CSR_PMPCFG2 = 12'h3A2;
	localparam [11:0] CSR_PMPCFG3 = 12'h3A3;
	localparam [11:0] CSR_PMPADDR0 = 12'h3B0;
	localparam [11:0] CSR_PMPADDR1 = 12'h3B1;
	localparam [11:0] CSR_PMPADDR2 = 12'h3B2;
	localparam [11:0] CSR_PMPADDR3 = 12'h3B3;
	localparam [11:0] CSR_PMPADDR4 = 12'h3B4;
	localparam [11:0] CSR_PMPADDR5 = 12'h3B5;
	localparam [11:0] CSR_PMPADDR6 = 12'h3B6;
	localparam [11:0] CSR_PMPADDR7 = 12'h3B7;
	localparam [11:0] CSR_PMPADDR8 = 12'h3B8;
	localparam [11:0] CSR_PMPADDR9 = 12'h3B9;
	localparam [11:0] CSR_PMPADDR10 = 12'h3BA;
	localparam [11:0] CSR_PMPADDR11 = 12'h3BB;
	localparam [11:0] CSR_PMPADDR12 = 12'h3BC;
	localparam [11:0] CSR_PMPADDR13 = 12'h3BD;
	localparam [11:0] CSR_PMPADDR14 = 12'h3BE;
	localparam [11:0] CSR_PMPADDR15 = 12'h3BF;
	localparam [11:0] CSR_DCSR = 12'h7b0;
	localparam [11:0] CSR_DPC = 12'h7b1;
	localparam [11:0] CSR_DSCRATCH0 = 12'h7b2;
	localparam [11:0] CSR_DSCRATCH1 = 12'h7b3;
	localparam [11:0] CSR_MCYCLE = 12'hB00;
	localparam [11:0] CSR_MINSTRET = 12'hB02;
	localparam [11:0] CSR_MCYCLEH = 12'hB80;
	localparam [11:0] CSR_MINSTRETH = 12'hB82;
	localparam [11:0] CSR_MHARTID = 12'hF14;
	localparam [4:0] ALU_GTU = 13;
	localparam [4:0] ALU_GE = 14;
	localparam [4:0] ALU_GEU = 15;
	localparam [4:0] ALU_EQ = 16;
	localparam [4:0] ALU_NE = 17;
	localparam [4:0] ALU_SLT = 18;
	localparam [4:0] ALU_SLTU = 19;
	localparam [1:0] CSR_OP_SET = 2;
	localparam [1:0] EXC_PC_DBD = 2;
	localparam [1:0] MD_OP_DIV = 2;
	localparam [1:0] OP_A_CURRPC = 2;
	localparam [1:0] RF_WD_CSR = 2;
	localparam [2:0] IMM_B_B = 2;
	localparam [2:0] PC_EXC = 2;
	localparam [4:0] ALU_XOR = 2;
	localparam [1:0] PMP_ACC_EXEC = 2'b00;
	localparam [1:0] PMP_MODE_OFF = 2'b00;
	localparam [1:0] PRIV_LVL_U = 2'b00;
	localparam [1:0] PMP_ACC_WRITE = 2'b01;
	localparam [1:0] PMP_MODE_TOR = 2'b01;
	localparam [1:0] PRIV_LVL_S = 2'b01;
	localparam [1:0] PMP_ACC_READ = 2'b10;
	localparam [1:0] PMP_MODE_NA4 = 2'b10;
	localparam [1:0] PRIV_LVL_H = 2'b10;
	localparam [1:0] PMP_MODE_NAPOT = 2'b11;
	localparam [1:0] PRIV_LVL_M = 2'b11;
	localparam [4:0] ALU_SLET = 20;
	localparam [4:0] ALU_SLETU = 21;
	localparam [1:0] CSR_OP_CLEAR = 3;
	localparam [1:0] EXC_PC_DBG_EXC = 3;
	localparam [1:0] MD_OP_REM = 3;
	localparam [1:0] OP_A_IMM = 3;
	localparam [2:0] IMM_B_U = 3;
	localparam [2:0] PC_ERET = 3;
	localparam [4:0] ALU_OR = 3;
	localparam [2:0] DBG_CAUSE_NONE = 3'h0;
	localparam [2:0] DBG_CAUSE_EBREAK = 3'h1;
	localparam [2:0] DBG_CAUSE_TRIGGER = 3'h2;
	localparam [2:0] DBG_CAUSE_HALTREQ = 3'h3;
	localparam [2:0] DBG_CAUSE_STEP = 3'h4;
	localparam [2:0] IMM_B_J = 4;
	localparam [2:0] PC_DRET = 4;
	localparam [4:0] ALU_AND = 4;
	localparam [3:0] XDEBUGVER_NO = 4'd0;
	localparam [3:0] XDEBUGVER_NONSTD = 4'd15;
	localparam [3:0] XDEBUGVER_STD = 4'd4;
	localparam [2:0] IMM_B_INCR_PC = 5;
	localparam [4:0] ALU_SRA = 5;
	localparam [2:0] IMM_B_INCR_ADDR = 6;
	localparam [4:0] ALU_SRL = 6;
	localparam [4:0] ALU_SLL = 7;
	localparam [6:0] OPCODE_LOAD = 7'h03;
	localparam [6:0] OPCODE_MISC_MEM = 7'h0f;
	localparam [6:0] OPCODE_OP_IMM = 7'h13;
	localparam [6:0] OPCODE_AUIPC = 7'h17;
	localparam [6:0] OPCODE_STORE = 7'h23;
	localparam [6:0] OPCODE_OP = 7'h33;
	localparam [6:0] OPCODE_LUI = 7'h37;
	localparam [6:0] OPCODE_BRANCH = 7'h63;
	localparam [6:0] OPCODE_JALR = 7'h67;
	localparam [6:0] OPCODE_JAL = 7'h6f;
	localparam [6:0] OPCODE_SYSTEM = 7'h73;
	localparam [4:0] ALU_LT = 8;
	localparam [4:0] ALU_LTU = 9;
	localparam [5:0] EXC_CAUSE_INSN_ADDR_MISA = {1'b0, 5'd00};
	localparam [5:0] EXC_CAUSE_INSTR_ACCESS_FAULT = {1'b0, 5'd01};
	localparam [5:0] EXC_CAUSE_ILLEGAL_INSN = {1'b0, 5'd02};
	localparam [5:0] EXC_CAUSE_BREAKPOINT = {1'b0, 5'd03};
	localparam [5:0] EXC_CAUSE_LOAD_ACCESS_FAULT = {1'b0, 5'd05};
	localparam [5:0] EXC_CAUSE_STORE_ACCESS_FAULT = {1'b0, 5'd07};
	localparam [5:0] EXC_CAUSE_ECALL_UMODE = {1'b0, 5'd08};
	localparam [5:0] EXC_CAUSE_ECALL_MMODE = {1'b0, 5'd11};
	localparam [5:0] EXC_CAUSE_IRQ_SOFTWARE_M = {1'b1, 5'd03};
	localparam [5:0] EXC_CAUSE_IRQ_TIMER_M = {1'b1, 5'd07};
	localparam [5:0] EXC_CAUSE_IRQ_EXTERNAL_M = {1'b1, 5'd11};
	localparam [5:0] EXC_CAUSE_IRQ_NM = {1'b1, 5'd31};
	localparam [1:0] MXL = 2'd1;
	localparam [31:0] MISA_VALUE = ((((((((((((0 << 0) | (1 << 2)) | (0 << 3)) | (sv2v_cast_32(RV32E) << 4)) | (0 << 5)) | (1 << 8)) | (sv2v_cast_32(RV32M) << 12)) | (0 << 13)) | (0 << 18)) | (0 << 20)) | (0 << 23)) | (sv2v_cast_32(MXL) << 30));
	reg [31:0] exception_pc;
	reg [1:0] priv_lvl_q;
	reg [1:0] priv_lvl_d;
	reg [5:0] mstatus_q;
	reg [5:0] mstatus_d;
	reg [17:0] mie_q;
	reg [17:0] mie_d;
	reg [31:0] mscratch_q;
	reg [31:0] mscratch_d;
	reg [31:0] mepc_q;
	reg [31:0] mepc_d;
	reg [5:0] mcause_q;
	reg [5:0] mcause_d;
	reg [31:0] mtval_q;
	reg [31:0] mtval_d;
	reg [31:0] mtvec_q;
	reg [31:0] mtvec_d;
	wire [17:0] mip;
	reg [31:0] dcsr_q;
	reg [31:0] dcsr_d;
	reg [31:0] depc_q;
	reg [31:0] depc_d;
	reg [31:0] dscratch0_q;
	reg [31:0] dscratch0_d;
	reg [31:0] dscratch1_q;
	reg [31:0] dscratch1_d;
	reg [2:0] mstack_q;
	reg [2:0] mstack_d;
	reg [31:0] mstack_epc_q;
	reg [31:0] mstack_epc_d;
	reg [5:0] mstack_cause_q;
	reg [5:0] mstack_cause_d;
	reg [31:0] pmp_addr_rdata [0:(PMP_MAX_REGIONS - 1)];
	wire [(PMP_CFG_W - 1):0] pmp_cfg_rdata [0:(PMP_MAX_REGIONS - 1)];
	reg [31:0] mcountinhibit_d;
	reg [31:0] mcountinhibit_q;
	wire [31:0] mcountinhibit;
	wire [31:0] mcountinhibit_force;
	reg mcountinhibit_we;
	reg [63:0] mhpmcounter_mask [0:(32 - 1)];
	reg [2047:0] mhpmcounter_d;
	reg [2047:0] mhpmcounter_q;
	reg [31:0] mhpmcounter_we;
	reg [31:0] mhpmcounterh_we;
	reg [31:0] mhpmcounter_incr;
	reg [31:0] mhpmevent [0:(32 - 1)];
	wire [4:0] mhpmcounter_idx;
	reg [31:0] csr_wdata_int;
	reg [31:0] csr_rdata_int;
	wire csr_we_int;
	reg csr_wreq;
	reg illegal_csr;
	wire illegal_csr_priv;
	wire illegal_csr_write;
	wire [7:0] unused_boot_addr;
	assign unused_boot_addr = boot_addr_i[7:0];
	wire [(12 - 1):0] csr_addr;
	assign csr_addr = csr_addr_i;
	assign mhpmcounter_idx = csr_addr[4:0];
	assign illegal_csr_priv = (csr_addr[9:8] > priv_lvl_q);
	assign illegal_csr_write = ((csr_addr[11:10] == 2'b11) && csr_wreq);
	assign illegal_csr_insn_o = (csr_access_i & ((illegal_csr | illegal_csr_write) | illegal_csr_priv));
	assign mip[17:17] = (irq_software_i & mie_q[17:17]);
	assign mip[16:16] = (irq_timer_i & mie_q[16:16]);
	assign mip[15:15] = (irq_external_i & mie_q[15:15]);
	assign mip[14:0] = (irq_fast_i & mie_q[14:0]);
	always @(*) begin
		csr_rdata_int = 1'sb0;
		illegal_csr = 1'b0;
		case (csr_addr_i)
			CSR_MHARTID: csr_rdata_int = hart_id_i;
			CSR_MSTATUS: begin
				csr_rdata_int = 1'sb0;
				csr_rdata_int[CSR_MSTATUS_MIE_BIT] = mstatus_q[5:5];
				csr_rdata_int[CSR_MSTATUS_MPIE_BIT] = mstatus_q[4:4];
				csr_rdata_int[CSR_MSTATUS_MPP_BIT_HIGH:CSR_MSTATUS_MPP_BIT_LOW] = mstatus_q[3:2];
				csr_rdata_int[CSR_MSTATUS_MPRV_BIT] = mstatus_q[1:1];
				csr_rdata_int[CSR_MSTATUS_TW_BIT] = mstatus_q[0:0];
			end
			CSR_MISA: csr_rdata_int = MISA_VALUE;
			CSR_MIE: begin
				csr_rdata_int = 1'sb0;
				csr_rdata_int[CSR_MSIX_BIT] = mie_q[17:17];
				csr_rdata_int[CSR_MTIX_BIT] = mie_q[16:16];
				csr_rdata_int[CSR_MEIX_BIT] = mie_q[15:15];
				csr_rdata_int[CSR_MFIX_BIT_HIGH:CSR_MFIX_BIT_LOW] = mie_q[14:0];
			end
			CSR_MSCRATCH: csr_rdata_int = mscratch_q;
			CSR_MTVEC: csr_rdata_int = mtvec_q;
			CSR_MEPC: csr_rdata_int = mepc_q;
			CSR_MCAUSE: csr_rdata_int = {mcause_q[5], 26'b0, mcause_q[4:0]};
			CSR_MTVAL: csr_rdata_int = mtval_q;
			CSR_MIP: begin
				csr_rdata_int = 1'sb0;
				csr_rdata_int[CSR_MSIX_BIT] = mip[17:17];
				csr_rdata_int[CSR_MTIX_BIT] = mip[16:16];
				csr_rdata_int[CSR_MEIX_BIT] = mip[15:15];
				csr_rdata_int[CSR_MFIX_BIT_HIGH:CSR_MFIX_BIT_LOW] = mip[14:0];
			end
			CSR_PMPCFG0: csr_rdata_int = {pmp_cfg_rdata[3], pmp_cfg_rdata[2], pmp_cfg_rdata[1], pmp_cfg_rdata[0]};
			CSR_PMPCFG1: csr_rdata_int = {pmp_cfg_rdata[7], pmp_cfg_rdata[6], pmp_cfg_rdata[5], pmp_cfg_rdata[4]};
			CSR_PMPCFG2: csr_rdata_int = {pmp_cfg_rdata[11], pmp_cfg_rdata[10], pmp_cfg_rdata[9], pmp_cfg_rdata[8]};
			CSR_PMPCFG3: csr_rdata_int = {pmp_cfg_rdata[15], pmp_cfg_rdata[14], pmp_cfg_rdata[13], pmp_cfg_rdata[12]};
			CSR_PMPADDR0: csr_rdata_int = pmp_addr_rdata[0];
			CSR_PMPADDR1: csr_rdata_int = pmp_addr_rdata[1];
			CSR_PMPADDR2: csr_rdata_int = pmp_addr_rdata[2];
			CSR_PMPADDR3: csr_rdata_int = pmp_addr_rdata[3];
			CSR_PMPADDR4: csr_rdata_int = pmp_addr_rdata[4];
			CSR_PMPADDR5: csr_rdata_int = pmp_addr_rdata[5];
			CSR_PMPADDR6: csr_rdata_int = pmp_addr_rdata[6];
			CSR_PMPADDR7: csr_rdata_int = pmp_addr_rdata[7];
			CSR_PMPADDR8: csr_rdata_int = pmp_addr_rdata[8];
			CSR_PMPADDR9: csr_rdata_int = pmp_addr_rdata[9];
			CSR_PMPADDR10: csr_rdata_int = pmp_addr_rdata[10];
			CSR_PMPADDR11: csr_rdata_int = pmp_addr_rdata[11];
			CSR_PMPADDR12: csr_rdata_int = pmp_addr_rdata[12];
			CSR_PMPADDR13: csr_rdata_int = pmp_addr_rdata[13];
			CSR_PMPADDR14: csr_rdata_int = pmp_addr_rdata[14];
			CSR_PMPADDR15: csr_rdata_int = pmp_addr_rdata[15];
			CSR_DCSR: begin
				csr_rdata_int = dcsr_q;
				illegal_csr = ~debug_mode_i;
			end
			CSR_DPC: begin
				csr_rdata_int = depc_q;
				illegal_csr = ~debug_mode_i;
			end
			CSR_DSCRATCH0: begin
				csr_rdata_int = dscratch0_q;
				illegal_csr = ~debug_mode_i;
			end
			CSR_DSCRATCH1: begin
				csr_rdata_int = dscratch1_q;
				illegal_csr = ~debug_mode_i;
			end
			CSR_MCOUNTINHIBIT: csr_rdata_int = mcountinhibit;
			CSR_MCYCLE: csr_rdata_int = mhpmcounter_q[1984+:32];
			CSR_MCYCLEH: csr_rdata_int = mhpmcounter_q[2016+:32];
			CSR_MINSTRET: csr_rdata_int = mhpmcounter_q[1856+:32];
			CSR_MINSTRETH: csr_rdata_int = mhpmcounter_q[1888+:32];
			default: if (((csr_addr & CSR_MASK_MCOUNTER) == CSR_OFF_MCOUNTER_SETUP)) begin
			csr_rdata_int = mhpmevent[mhpmcounter_idx];
			if ((((csr_addr[4:0] == 5'b00000) || (csr_addr[4:0] == 5'b00001)) || (csr_addr[4:0] == 5'b00010)))
				illegal_csr = 1'b1;
		end
		else if (((csr_addr & CSR_MASK_MCOUNTER) == CSR_OFF_MCOUNTER)) begin
			csr_rdata_int = mhpmcounter_q[((31 - mhpmcounter_idx) * 64)+:32];
			if ((((csr_addr[4:0] == 5'b00000) || (csr_addr[4:0] == 5'b00001)) || (csr_addr[4:0] == 5'b00010)))
				illegal_csr = 1'b1;
		end
		else if (((csr_addr & CSR_MASK_MCOUNTER) == CSR_OFF_MCOUNTERH)) begin
			csr_rdata_int = mhpmcounter_q[(((31 - mhpmcounter_idx) * 64) + 32)+:32];
			if ((((csr_addr[4:0] == 5'b00000) || (csr_addr[4:0] == 5'b00001)) || (csr_addr[4:0] == 5'b00010)))
				illegal_csr = 1'b1;
		end
		else
			illegal_csr = 1'b1;
		endcase
	end
	always @(*) begin
		exception_pc = pc_id_i;
		priv_lvl_d = priv_lvl_q;
		mstatus_d = mstatus_q;
		mie_d = mie_q;
		mscratch_d = mscratch_q;
		mepc_d = mepc_q;
		mcause_d = mcause_q;
		mtval_d = mtval_q;
		mtvec_d = (csr_mtvec_init_i ? {boot_addr_i[31:8], 6'b0, 2'b01} : mtvec_q);
		dcsr_d = dcsr_q;
		depc_d = depc_q;
		dscratch0_d = dscratch0_q;
		dscratch1_d = dscratch1_q;
		mstack_d = mstack_q;
		mstack_epc_d = mstack_epc_q;
		mstack_cause_d = mstack_cause_q;
		mcountinhibit_we = 1'b0;
		mhpmcounter_we = 1'sb0;
		mhpmcounterh_we = 1'sb0;
		if (csr_we_int)
			case (csr_addr_i)
				CSR_MSTATUS: begin
					mstatus_d = sv2v_struct_BF3E9(csr_wdata_int[CSR_MSTATUS_MIE_BIT], csr_wdata_int[CSR_MSTATUS_MPIE_BIT], csr_wdata_int[CSR_MSTATUS_MPP_BIT_HIGH:CSR_MSTATUS_MPP_BIT_LOW], csr_wdata_int[CSR_MSTATUS_MPRV_BIT], csr_wdata_int[CSR_MSTATUS_TW_BIT]);
					if (((mstatus_d[3:2] != PRIV_LVL_M) && (mstatus_d[3:2] != PRIV_LVL_U)))
						mstatus_d[3:2] = PRIV_LVL_M;
				end
				CSR_MIE: begin
					mie_d[17:17] = csr_wdata_int[CSR_MSIX_BIT];
					mie_d[16:16] = csr_wdata_int[CSR_MTIX_BIT];
					mie_d[15:15] = csr_wdata_int[CSR_MEIX_BIT];
					mie_d[14:0] = csr_wdata_int[CSR_MFIX_BIT_HIGH:CSR_MFIX_BIT_LOW];
				end
				CSR_MSCRATCH: mscratch_d = csr_wdata_int;
				CSR_MEPC: mepc_d = {csr_wdata_int[31:1], 1'b0};
				CSR_MCAUSE: mcause_d = {csr_wdata_int[31], csr_wdata_int[4:0]};
				CSR_MTVAL: mtval_d = csr_wdata_int;
				CSR_MTVEC: mtvec_d = {csr_wdata_int[31:8], 6'b0, 2'b01};
				CSR_DCSR: begin
					dcsr_d = csr_wdata_int;
					dcsr_d[31:28] = XDEBUGVER_STD;
					if (((dcsr_d[1:0] != PRIV_LVL_M) && (dcsr_d[1:0] != PRIV_LVL_U)))
						dcsr_d[1:0] = PRIV_LVL_M;
					dcsr_d[3:3] = 1'b0;
					dcsr_d[4:4] = 1'b0;
					dcsr_d[10:10] = 1'b0;
					dcsr_d[9:9] = 1'b0;
					dcsr_d[5:5] = 1'b0;
					dcsr_d[14:14] = 1'b0;
					dcsr_d[27:16] = 12'h0;
				end
				CSR_DPC:
					if ((csr_wdata_int[0] == 1'b0))
						depc_d = csr_wdata_int;
				CSR_DSCRATCH0: dscratch0_d = csr_wdata_int;
				CSR_DSCRATCH1: dscratch1_d = csr_wdata_int;
				CSR_MCOUNTINHIBIT: mcountinhibit_we = 1'b1;
				CSR_MCYCLE: mhpmcounter_we[0] = 1'b1;
				CSR_MCYCLEH: mhpmcounterh_we[0] = 1'b1;
				CSR_MINSTRET: mhpmcounter_we[2] = 1'b1;
				CSR_MINSTRETH: mhpmcounterh_we[2] = 1'b1;
				default: if (((csr_addr & CSR_MASK_MCOUNTER) == CSR_OFF_MCOUNTER))
				mhpmcounter_we[mhpmcounter_idx] = 1'b1;
			else if (((csr_addr & CSR_MASK_MCOUNTER) == CSR_OFF_MCOUNTERH))
				mhpmcounterh_we[mhpmcounter_idx] = 1'b1;
			endcase
		case (1'b1)
			csr_save_cause_i: begin
				case (1'b1)
					csr_save_if_i: exception_pc = pc_if_i;
					csr_save_id_i: exception_pc = pc_id_i;
					default: ;
				endcase
				if (debug_csr_save_i) begin
					dcsr_d[1:0] = priv_lvl_q;
					dcsr_d[8:6] = debug_cause_i;
					depc_d = exception_pc;
				end
				else begin
					priv_lvl_d = PRIV_LVL_M;
					mtval_d = csr_mtval_i;
					mstatus_d[5:5] = 1'b0;
					mstatus_d[4:4] = mstatus_q[5:5];
					mstatus_d[3:2] = priv_lvl_q;
					mepc_d = exception_pc;
					mcause_d = csr_mcause_i;
					mstack_d[2:2] = mstatus_q[4:4];
					mstack_d[1:0] = mstatus_q[3:2];
					mstack_epc_d = mepc_q;
					mstack_cause_d = mcause_q;
				end
			end
			csr_restore_mret_i: begin
				priv_lvl_d = mstatus_q[3:2];
				mstatus_d[5:5] = mstatus_q[4:4];
				mstatus_d[4:4] = mstack_q[2:2];
				mstatus_d[3:2] = mstack_q[1:0];
				mepc_d = mstack_epc_q;
				mcause_d = mstack_cause_q;
				mstack_d[2:2] = 1'b1;
				mstack_d[1:0] = PRIV_LVL_U;
			end
			default: ;
		endcase
	end
	always @(*) begin
		csr_wreq = 1'b1;
		case (csr_op_i)
			CSR_OP_WRITE: csr_wdata_int = csr_wdata_i;
			CSR_OP_SET: csr_wdata_int = (csr_wdata_i | csr_rdata_o);
			CSR_OP_CLEAR: csr_wdata_int = (~csr_wdata_i & csr_rdata_o);
			CSR_OP_READ: begin
				csr_wdata_int = csr_wdata_i;
				csr_wreq = 1'b0;
			end
			default: begin
			csr_wdata_int = 1'sbX;
			csr_wreq = 1'bX;
		end
		endcase
	end
	assign csr_we_int = ((csr_wreq & ~illegal_csr_insn_o) & instr_new_id_i);
	assign csr_rdata_o = csr_rdata_int;
	assign csr_msip_o = mip[17:17];
	assign csr_mtip_o = mip[16:16];
	assign csr_meip_o = mip[15:15];
	assign csr_mfip_o = mip[14:0];
	assign csr_mepc_o = mepc_q;
	assign csr_depc_o = depc_q;
	assign csr_mtvec_o = mtvec_q;
	assign csr_mstatus_mie_o = mstatus_q[5:5];
	assign csr_mstatus_tw_o = mstatus_q[0:0];
	assign debug_single_step_o = dcsr_q[2:2];
	assign debug_ebreakm_o = dcsr_q[15:15];
	assign debug_ebreaku_o = dcsr_q[12:12];
	assign irq_pending_o = (((csr_msip_o | csr_mtip_o) | csr_meip_o) | |csr_mfip_o);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			priv_lvl_q <= PRIV_LVL_M;
			mstatus_q <= sv2v_struct_BF3E9(1'b0, 1'b1, PRIV_LVL_U, 1'b0, 1'b0);
			mie_q <= 1'sb0;
			mscratch_q <= 1'sb0;
			mepc_q <= 1'sb0;
			mcause_q <= 1'sb0;
			mtval_q <= 1'sb0;
			mtvec_q <= 32'b01;
			dcsr_q <= sv2v_struct_996E9(XDEBUGVER_STD, 1'sb0, 1'sb0, 1'sb0, 1'sb0, 1'sb0, 1'sb0, 1'sb0, 1'sb0, DBG_CAUSE_NONE, 1'sb0, 1'sb0, 1'sb0, 1'sb0, PRIV_LVL_M);
			depc_q <= 1'sb0;
			dscratch0_q <= 1'sb0;
			dscratch1_q <= 1'sb0;
			mstack_q <= sv2v_struct_70E1D(1'b1, PRIV_LVL_U);
			mstack_epc_q <= 1'sb0;
			mstack_cause_q <= 1'sb0;
		end
		else begin
			priv_lvl_q <= priv_lvl_d;
			mstatus_q <= mstatus_d;
			mie_q <= mie_d;
			mscratch_q <= mscratch_d;
			mepc_q <= mepc_d;
			mcause_q <= mcause_d;
			mtval_q <= mtval_d;
			mtvec_q <= mtvec_d;
			dcsr_q <= dcsr_d;
			depc_q <= depc_d;
			dscratch0_q <= dscratch0_d;
			dscratch1_q <= dscratch1_d;
			mstack_q <= mstack_d;
			mstack_epc_q <= mstack_epc_d;
			mstack_cause_q <= mstack_cause_d;
		end
	assign priv_mode_id_o = priv_lvl_q;
	assign priv_mode_if_o = priv_lvl_d;
	assign priv_mode_lsu_o = (mstatus_q[1:1] ? mstatus_q[3:2] : priv_lvl_q);
	generate
		if (PMPEnable) begin : g_pmp_registers
			reg [5:0] pmp_cfg [0:(PMPNumRegions - 1)];
			reg [5:0] pmp_cfg_wdata [0:(PMPNumRegions - 1)];
			reg [31:0] pmp_addr [0:(PMPNumRegions - 1)];
			wire [(PMPNumRegions - 1):0] pmp_cfg_we;
			wire [(PMPNumRegions - 1):0] pmp_addr_we;
			genvar g_exp_rd_data_i;
			for (g_exp_rd_data_i = 0; (g_exp_rd_data_i < PMP_MAX_REGIONS); g_exp_rd_data_i = (g_exp_rd_data_i + 1)) begin : g_exp_rd_data
				if ((g_exp_rd_data_i < PMPNumRegions)) begin : g_implemented_regions
					assign pmp_cfg_rdata[g_exp_rd_data_i] = {pmp_cfg[g_exp_rd_data_i][5:5], 2'b00, pmp_cfg[g_exp_rd_data_i][4:3], pmp_cfg[g_exp_rd_data_i][2:2], pmp_cfg[g_exp_rd_data_i][1:1], pmp_cfg[g_exp_rd_data_i][0:0]};
					if ((PMPGranularity == 0)) begin : g_pmp_g0
						always @(*) pmp_addr_rdata[g_exp_rd_data_i] = pmp_addr[g_exp_rd_data_i];
					end
					else if ((PMPGranularity == 1)) begin : g_pmp_g1
						always @(*) begin
							pmp_addr_rdata[g_exp_rd_data_i] = pmp_addr[g_exp_rd_data_i];
							if (((pmp_cfg[g_exp_rd_data_i][4:3] == PMP_MODE_OFF) || (pmp_cfg[g_exp_rd_data_i][4:3] == PMP_MODE_TOR)))
								pmp_addr_rdata[g_exp_rd_data_i][(PMPGranularity - 1):0] = 1'sb0;
						end
					end
					else begin : g_pmp_g2
						always @(*) begin
							pmp_addr_rdata[g_exp_rd_data_i] = pmp_addr[g_exp_rd_data_i];
							if (((pmp_cfg[g_exp_rd_data_i][4:3] == PMP_MODE_OFF) || (pmp_cfg[g_exp_rd_data_i][4:3] == PMP_MODE_TOR)))
								pmp_addr_rdata[g_exp_rd_data_i][(PMPGranularity - 1):0] = 1'sb0;
							else if ((pmp_cfg[g_exp_rd_data_i][4:3] == PMP_MODE_NAPOT))
								pmp_addr_rdata[g_exp_rd_data_i][(PMPGranularity - 2):0] = 1'sb1;
						end
					end
				end
				else begin : g_other_regions
					assign pmp_cfg_rdata[g_exp_rd_data_i] = 1'sb0;
					always @(*) pmp_addr_rdata[g_exp_rd_data_i] = 1'sb0;
				end
			end
			genvar g_pmp_csrs_i;
			for (g_pmp_csrs_i = 0; (g_pmp_csrs_i < PMPNumRegions); g_pmp_csrs_i = (g_pmp_csrs_i + 1)) begin : g_pmp_csrs
				assign pmp_cfg_we[g_pmp_csrs_i] = ((csr_we_int & ~pmp_cfg[g_pmp_csrs_i][5:5]) & (csr_addr == (CSR_OFF_PMP_CFG + (g_pmp_csrs_i[11:0] >> 2))));
				always @(*) pmp_cfg_wdata[g_pmp_csrs_i][5:5] = csr_wdata_int[(((g_pmp_csrs_i % 4) * PMP_CFG_W) + 7)];
				always @(*)
					case (csr_wdata_int[(((g_pmp_csrs_i % 4) * PMP_CFG_W) + 3)+:2])
						2'b00: pmp_cfg_wdata[g_pmp_csrs_i][4:3] = PMP_MODE_OFF;
						2'b01: pmp_cfg_wdata[g_pmp_csrs_i][4:3] = PMP_MODE_TOR;
						2'b10: pmp_cfg_wdata[g_pmp_csrs_i][4:3] = ((PMPGranularity == 0) ? PMP_MODE_NA4 : PMP_MODE_OFF);
						2'b11: pmp_cfg_wdata[g_pmp_csrs_i][4:3] = PMP_MODE_NAPOT;
						default: pmp_cfg_wdata[g_pmp_csrs_i][4:3] = 1'sbX;
					endcase
				always @(*) pmp_cfg_wdata[g_pmp_csrs_i][2:2] = csr_wdata_int[(((g_pmp_csrs_i % 4) * PMP_CFG_W) + 2)];
				always @(*) pmp_cfg_wdata[g_pmp_csrs_i][1:1] = &csr_wdata_int[((g_pmp_csrs_i % 4) * PMP_CFG_W)+:2];
				always @(*) pmp_cfg_wdata[g_pmp_csrs_i][0:0] = csr_wdata_int[((g_pmp_csrs_i % 4) * PMP_CFG_W)];
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni)
						pmp_cfg[g_pmp_csrs_i] <= 'b0;
					else if (pmp_cfg_we[g_pmp_csrs_i])
						pmp_cfg[g_pmp_csrs_i] <= pmp_cfg_wdata[g_pmp_csrs_i];
				if ((g_pmp_csrs_i < (PMPNumRegions - 1))) begin : g_lower
					assign pmp_addr_we[g_pmp_csrs_i] = (((csr_we_int & ~pmp_cfg[g_pmp_csrs_i][5:5]) & (pmp_cfg[(g_pmp_csrs_i + 1)][4:3] != PMP_MODE_TOR)) & (csr_addr == (CSR_OFF_PMP_ADDR + g_pmp_csrs_i[11:0])));
				end
				else begin : g_upper
					assign pmp_addr_we[g_pmp_csrs_i] = ((csr_we_int & ~pmp_cfg[g_pmp_csrs_i][5:5]) & (csr_addr == (CSR_OFF_PMP_ADDR + g_pmp_csrs_i[11:0])));
				end
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni)
						pmp_addr[g_pmp_csrs_i] <= 'b0;
					else if (pmp_addr_we[g_pmp_csrs_i])
						pmp_addr[g_pmp_csrs_i] <= csr_wdata_int;
				assign csr_pmp_cfg_o[(((0 >= (PMPNumRegions - 1)) ? g_pmp_csrs_i : ((PMPNumRegions - 1) - g_pmp_csrs_i)) * 6)+:6] = pmp_cfg[g_pmp_csrs_i];
				assign csr_pmp_addr_o[(((0 >= (PMPNumRegions - 1)) ? g_pmp_csrs_i : ((PMPNumRegions - 1) - g_pmp_csrs_i)) * 34)+:34] = {pmp_addr[g_pmp_csrs_i], 2'b00};
			end
		end
		else begin : g_no_pmp_tieoffs
			genvar g_rdata_i;
			for (g_rdata_i = 0; (g_rdata_i < PMP_MAX_REGIONS); g_rdata_i = (g_rdata_i + 1)) begin : g_rdata
				always @(*) pmp_addr_rdata[g_rdata_i] = 1'sb0;
				assign pmp_cfg_rdata[g_rdata_i] = 1'sb0;
			end
			genvar g_outputs_i;
			for (g_outputs_i = 0; (g_outputs_i < PMPNumRegions); g_outputs_i = (g_outputs_i + 1)) begin : g_outputs
				assign csr_pmp_cfg_o[(((0 >= (PMPNumRegions - 1)) ? g_outputs_i : ((PMPNumRegions - 1) - g_outputs_i)) * 6)+:6] = 1'b0;
				assign csr_pmp_addr_o[(((0 >= (PMPNumRegions - 1)) ? g_outputs_i : ((PMPNumRegions - 1) - g_outputs_i)) * 34)+:34] = 1'sb0;
			end
		end
	endgenerate
	always @(*) begin : mcountinhibit_update
		if ((mcountinhibit_we == 1'b1))
			mcountinhibit_d = {csr_wdata_int[31:2], 1'b0, csr_wdata_int[0]};
		else
			mcountinhibit_d = mcountinhibit_q;
	end
	assign mcountinhibit_force = {{(29 - MHPMCounterNum) {1'b1}}, {MHPMCounterNum {1'b0}}, 3'b000};
	assign mcountinhibit = (mcountinhibit_q | mcountinhibit_force);
	always @(*) begin : gen_mhpmcounter_incr
		mhpmcounter_incr[0] = 1'b1;
		mhpmcounter_incr[1] = 1'b0;
		mhpmcounter_incr[2] = instr_ret_i;
		mhpmcounter_incr[3] = lsu_busy_i;
		mhpmcounter_incr[4] = (imiss_i & ~pc_set_i);
		mhpmcounter_incr[5] = mem_load_i;
		mhpmcounter_incr[6] = mem_store_i;
		mhpmcounter_incr[7] = jump_i;
		mhpmcounter_incr[8] = branch_i;
		mhpmcounter_incr[9] = branch_taken_i;
		mhpmcounter_incr[10] = instr_ret_compressed_i;
		begin : sv2v_autoblock_14
			reg [31:0] i;
			for (i = (3 + MHPMCounterNum); (i < 32); i = (i + 1))
				begin : gen_mhpmcounter_incr_inactive
					mhpmcounter_incr[i] = 1'b0;
				end
		end
	end
	always @(*) begin : gen_mhpmevent
		begin : sv2v_autoblock_15
			reg signed [31:0] i;
			for (i = 0; (i < 32); i = (i + 1))
				begin : gen_mhpmevent_active
					mhpmevent[i] = 1'sb0;
					mhpmevent[i][i] = 1'b1;
				end
		end
		mhpmevent[1] = 1'sb0;
		begin : sv2v_autoblock_16
			reg [31:0] i;
			for (i = (3 + MHPMCounterNum); (i < 32); i = (i + 1))
				begin : gen_mhpmevent_inactive
					mhpmevent[i] = 1'sb0;
				end
		end
	end
	always @(*) begin : gen_mask
		begin : sv2v_autoblock_17
			reg signed [31:0] i;
			for (i = 0; (i < 3); i = (i + 1))
				begin : gen_mask_fixed
					mhpmcounter_mask[i] = {64 {1'b1}};
				end
		end
		begin : sv2v_autoblock_18
			reg [31:0] i;
			for (i = 3; (i < (3 + MHPMCounterNum)); i = (i + 1))
				begin : gen_mask_configurable
					mhpmcounter_mask[i] = {{(64 - MHPMCounterWidth) {1'b0}}, {MHPMCounterWidth {1'b1}}};
				end
		end
		begin : sv2v_autoblock_19
			reg [31:0] i;
			for (i = (3 + MHPMCounterNum); (i < 32); i = (i + 1))
				begin : gen_mask_inactive
					mhpmcounter_mask[i] = 1'sb0;
				end
		end
	end
	always @(*) begin : mhpmcounter_update
		mhpmcounter_d = mhpmcounter_q;
		begin : sv2v_autoblock_20
			reg signed [31:0] i;
			for (i = 0; (i < 32); i = (i + 1))
				begin : gen_mhpmcounter_update
					if ((mhpmcounter_incr[i] & ~mcountinhibit[i]))
						mhpmcounter_d[((31 - i) * 64)+:64] = (mhpmcounter_mask[i] & (mhpmcounter_q[((31 - i) * 64)+:64] + 64'h1));
					if (mhpmcounter_we[i])
						mhpmcounter_d[((31 - i) * 64)+:32] = (mhpmcounter_mask[i][31:0] & csr_wdata_int);
					else if (mhpmcounterh_we[i])
						mhpmcounter_d[(((31 - i) * 64) + 32)+:32] = (mhpmcounter_mask[i][63:32] & csr_wdata_int);
				end
		end
	end
	always @(posedge clk_i or negedge rst_ni) begin : perf_counter_registers
		if (!rst_ni) begin
			mcountinhibit_q <= 1'sb0;
			begin : sv2v_autoblock_21
				reg signed [31:0] i;
				for (i = 0; (i < 32); i = (i + 1))
					mhpmcounter_q[((31 - i) * 64)+:64] <= 1'sb0;
			end
		end
		else begin
			mhpmcounter_q <= mhpmcounter_d;
			mcountinhibit_q <= mcountinhibit_d;
		end
	end
	function [5:0] sv2v_struct_BF3E9;
		input reg mie;
		input reg mpie;
		input reg [1:0] mpp;
		input reg mprv;
		input reg tw;
		sv2v_struct_BF3E9 = {mie, mpie, mpp, mprv, tw};
	endfunction
	function [2:0] sv2v_struct_70E1D;
		input reg mpie;
		input reg [1:0] mpp;
		sv2v_struct_70E1D = {mpie, mpp};
	endfunction
	function [31:0] sv2v_struct_996E9;
		input reg [3:0] xdebugver;
		input reg [11:0] zero2;
		input reg ebreakm;
		input reg zero1;
		input reg ebreaks;
		input reg ebreaku;
		input reg stepie;
		input reg stopcount;
		input reg stoptime;
		input reg [2:0] cause;
		input reg zero0;
		input reg mprven;
		input reg nmip;
		input reg step;
		input reg [1:0] prv;
		sv2v_struct_996E9 = {xdebugver, zero2, ebreakm, zero1, ebreaks, ebreaku, stepie, stopcount, stoptime, cause, zero0, mprven, nmip, step, prv};
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
endmodule

module usbuart_usbif (
	clk_48mhz_i,
	rst_ni,
	usb_dp_o,
	usb_dn_o,
	usb_dp_i,
	usb_dn_i,
	usb_tx_en_o,
	tx_empty,
	rx_full,
	tx_read,
	rx_write,
	rx_err,
	rx_fifo_wdata,
	tx_fifo_rdata,
	rx_fifo_wdepth,
	status_frame_o,
	status_host_lost_o,
	status_host_timeout_o,
	status_device_address_o,
	parity_o,
	baud_o
);
	input clk_48mhz_i;
	input rst_ni;
	output usb_dp_o;
	output usb_dn_o;
	input usb_dp_i;
	input usb_dn_i;
	output usb_tx_en_o;
	input tx_empty;
	input rx_full;
	output tx_read;
	output rx_write;
	output rx_err;
	output [7:0] rx_fifo_wdata;
	input [7:0] tx_fifo_rdata;
	input [5:0] rx_fifo_wdepth;
	output reg [10:0] status_frame_o;
	output wire status_host_lost_o;
	output reg status_host_timeout_o;
	output wire [6:0] status_device_address_o;
	output wire [1:0] parity_o;
	output wire [15:0] baud_o;
	localparam MaxPktSizeByte = 32;
	localparam PktW = 5;
	localparam CtrlEp = 0;
	localparam FifoEp = 1;
	reg [5:0] ns_cnt;
	wire us_tick;
	assign us_tick = (ns_cnt == 6'd48);
	always @(posedge clk_48mhz_i or negedge rst_ni)
		if (!rst_ni)
			ns_cnt <= 1'sb0;
		else if (us_tick)
			ns_cnt <= 1'sb0;
		else
			ns_cnt <= (ns_cnt + 1'b1);
	wire [6:0] dev_addr;
	wire [7:0] out_ep_data;
	wire [3:0] in_ep_current;
	wire in_ep_rollback;
	wire in_ep_acked;
	wire [(PktW - 1):0] in_ep_get_addr;
	wire in_ep_data_get;
	wire [3:0] out_ep_current;
	wire out_ep_rollback;
	wire out_ep_acked;
	wire [(PktW - 1):0] out_ep_put_addr;
	wire out_ep_data_put;
	wire ctrl_out_ep_setup;
	wire ctrl_out_ep_stall;
	wire ctrl_out_ep_full;
	wire [7:0] ctrl_in_ep_data;
	wire ctrl_in_ep_data_done;
	wire ctrl_in_ep_stall;
	wire ctrl_in_ep_has_data;
	wire serial_out_ep_setup;
	wire serial_out_ep_stall;
	wire serial_out_ep_full;
	wire [7:0] serial_in_ep_data;
	wire serial_in_ep_data_done;
	wire serial_in_ep_stall;
	wire serial_in_ep_has_data;
	wire sof_valid;
	wire [10:0] frame_index_raw;
	reg [19:0] host_presence_timer;
	assign status_device_address_o = dev_addr;
	wire out_ctrl_put;
	wire out_ctrl_acked;
	wire out_ctrl_rollback;
	wire in_ctrl_get;
	wire in_ctrl_acked;
	wire in_ctrl_rollback;
	assign out_ctrl_put = (out_ep_data_put && (out_ep_current == CtrlEp));
	assign out_ctrl_acked = (out_ep_acked && (out_ep_current == CtrlEp));
	assign out_ctrl_rollback = (out_ep_rollback && (out_ep_current == CtrlEp));
	assign in_ctrl_get = (in_ep_data_get && (in_ep_current == CtrlEp));
	assign in_ctrl_acked = (in_ep_acked && (in_ep_current == CtrlEp));
	assign in_ctrl_rollback = (in_ep_rollback && (in_ep_current == CtrlEp));
	usb_serial_ctrl_ep #(.MaxPktSizeByte(MaxPktSizeByte)) u_usb_serial_ctrl_ep(
		.clk_i(clk_48mhz_i),
		.rst_ni(rst_ni),
		.dev_addr(dev_addr),
		.out_ep_data_put_i(out_ctrl_put),
		.out_ep_put_addr_i(out_ep_put_addr),
		.out_ep_data_i(out_ep_data),
		.out_ep_acked_i(out_ctrl_acked),
		.out_ep_rollback_i(out_ctrl_rollback),
		.out_ep_setup_i(ctrl_out_ep_setup),
		.out_ep_full_o(ctrl_out_ep_full),
		.out_ep_stall_o(ctrl_out_ep_stall),
		.in_ep_rollback_i(in_ctrl_rollback),
		.in_ep_acked_i(in_ctrl_acked),
		.in_ep_get_addr_i(in_ep_get_addr),
		.in_ep_data_get_i(in_ctrl_get),
		.in_ep_stall_o(ctrl_in_ep_stall),
		.in_ep_has_data_o(ctrl_in_ep_has_data),
		.in_ep_data_o(ctrl_in_ep_data[7:0]),
		.in_ep_data_done_o(ctrl_in_ep_data_done)
	);
	wire out_fifo_put;
	wire out_fifo_acked;
	wire out_fifo_rollback;
	wire in_fifo_get;
	wire in_fifo_acked;
	wire in_fifo_rollback;
	assign out_fifo_put = (out_ep_data_put && (out_ep_current == FifoEp));
	assign out_fifo_acked = (out_ep_acked && (out_ep_current == FifoEp));
	assign out_fifo_rollback = (out_ep_rollback && (out_ep_current == FifoEp));
	assign in_fifo_get = (in_ep_data_get && (in_ep_current == FifoEp));
	assign in_fifo_acked = (in_ep_acked && (in_ep_current == FifoEp));
	assign in_fifo_rollback = (in_ep_rollback && (in_ep_current == FifoEp));
	usb_serial_fifo_ep #(.MaxPktSizeByte(MaxPktSizeByte)) u_usb_serial_fifo_ep(
		.clk_i(clk_48mhz_i),
		.rst_ni(rst_ni),
		.out_ep_data_put_i(out_fifo_put),
		.out_ep_put_addr_i(out_ep_put_addr),
		.out_ep_data_i(out_ep_data),
		.out_ep_acked_i(out_fifo_acked),
		.out_ep_rollback_i(out_fifo_rollback),
		.out_ep_setup_i(serial_out_ep_setup),
		.out_ep_full_o(serial_out_ep_full),
		.out_ep_stall_o(serial_out_ep_stall),
		.in_ep_rollback_i(in_fifo_rollback),
		.in_ep_acked_i(in_fifo_acked),
		.in_ep_get_addr_i(in_ep_get_addr),
		.in_ep_data_get_i(in_fifo_get),
		.in_ep_stall_o(serial_in_ep_stall),
		.in_ep_has_data_o(serial_in_ep_has_data),
		.in_ep_data_o(serial_in_ep_data[7:0]),
		.in_ep_data_done_o(serial_in_ep_data_done),
		.tx_empty(tx_empty),
		.rx_full(rx_full),
		.tx_read(tx_read),
		.rx_write(rx_write),
		.rx_err(rx_err),
		.rx_fifo_wdata(rx_fifo_wdata),
		.tx_fifo_rdata(tx_fifo_rdata),
		.parity_o(parity_o),
		.baud_o(baud_o)
	);
	usb_fs_nb_pe #(
		.NumOutEps(2),
		.NumInEps(2),
		.MaxPktSizeByte(MaxPktSizeByte)
	) u_usb_fs_nb_pe(
		.clk_48mhz_i(clk_48mhz_i),
		.rst_ni(rst_ni),
		.link_reset_i(1'b0),
		.usb_p_tx_o(usb_dp_o),
		.usb_n_tx_o(usb_dn_o),
		.usb_p_rx_i(usb_dp_i),
		.usb_n_rx_i(usb_dn_i),
		.usb_tx_en_o(usb_tx_en_o),
		.dev_addr_i(dev_addr),
		.out_ep_current_o(out_ep_current),
		.out_ep_data_put_o(out_ep_data_put),
		.out_ep_put_addr_o(out_ep_put_addr),
		.out_ep_data_o(out_ep_data),
		.out_ep_acked_o(out_ep_acked),
		.out_ep_rollback_o(out_ep_rollback),
		.out_ep_newpkt_o(),
		.out_ep_setup_o({serial_out_ep_setup, ctrl_out_ep_setup}),
		.out_ep_full_i({serial_out_ep_full, ctrl_out_ep_full}),
		.out_ep_stall_i({serial_out_ep_stall, ctrl_out_ep_stall}),
		.in_ep_current_o(in_ep_current),
		.in_ep_rollback_o(in_ep_rollback),
		.in_ep_acked_o(in_ep_acked),
		.in_ep_get_addr_o(in_ep_get_addr),
		.in_ep_data_get_o(in_ep_data_get),
		.in_ep_newpkt_o(),
		.in_ep_stall_i({serial_in_ep_stall, ctrl_in_ep_stall}),
		.in_ep_has_data_i({serial_in_ep_has_data, ctrl_in_ep_has_data}),
		.in_ep_data_i(((in_ep_current == 4'b1) ? serial_in_ep_data : ctrl_in_ep_data)),
		.in_ep_data_done_i({serial_in_ep_data_done, ctrl_in_ep_data_done}),
		.sof_valid_o(sof_valid),
		.frame_index_o(frame_index_raw)
	);
	assign status_host_lost_o = (host_presence_timer[19:12] != 0);
	always @(posedge clk_48mhz_i or negedge rst_ni)
		if (!rst_ni) begin
			host_presence_timer <= 1'sb0;
			status_host_timeout_o <= 1'b0;
			status_frame_o <= 1'sb0;
		end
		else if (sof_valid) begin
			host_presence_timer <= 0;
			status_host_timeout_o <= 0;
			status_frame_o <= frame_index_raw;
		end
		else if ((host_presence_timer > 1000000))
			status_host_timeout_o <= 1;
		else if (us_tick)
			host_presence_timer <= (host_presence_timer + 1);
endmodule
